`timescale 1ns/1ps

module tb_commit_rename;

  // -------------------------
  // Parameters (match DUT)
  // -------------------------
  localparam int ARCH_REGS = 32;
  localparam int PHYS_REGS = 64;
  localparam int PHYS_W    = $clog2(PHYS_REGS);
  localparam int ROB_SIZE  = 16;
  localparam int ROB_W     = $clog2(ROB_SIZE);

  // -------------------------
  // Clock / Reset
  // -------------------------
  logic clk, rst_n;
  initial clk = 1'b0;
  always #5 clk = ~clk; // 100MHz

  // -------------------------
  // DUT I/O
  // -------------------------
  logic               alloc_valid;
  logic               alloc_ready;
  logic               alloc_uses_rd;
  logic [4:0]         alloc_rd_arch;
  logic               alloc_is_branch, alloc_is_load, alloc_is_store;
  logic [31:0]        alloc_pc;
  logic               alloc_epoch;
  logic [ROB_W-1:0]   alloc_rob_idx;

  logic               wb_valid;
  logic [ROB_W-1:0]   wb_rob_idx;
  logic               wb_epoch;

  logic               commit_valid;
  logic               commit_ready;

  logic               commit_uses_rd;
  logic [4:0]         commit_rd_arch;
  logic [PHYS_W-1:0]  commit_pd_new;
  logic [PHYS_W-1:0]  commit_pd_old;
  logic               commit_is_branch, commit_is_load, commit_is_store;

  logic               flush_valid;
  logic [ROB_W-1:0]   flush_rob_idx;
  logic               flush_epoch;

  logic [4:0]         rs1_arch, rs2_arch;

  // debug outputs from DUT (your file declares [4:0] widths; we cast to PHYS_W)
  wire  [PHYS_W-1:0]         rs1_phys_dbg;
  wire  [PHYS_W-1:0]         rs2_phys_dbg;
  wire  [PHYS_W-1:0]         rd_phys_dbg;
  wire  [PHYS_W-1:0]         rd_new_phys_dbg;

  // Cast to full phys width (safe for PHYS_REGS<=32? here PHYS_REGS=64 so debug is too narrow)
  // If your debug ports are truly 5 bits, they cannot represent 32..63. You should widen them to [PHYS_W-1:0].
  // For now we still cast; TB will warn if it sees truncation.
  logic [PHYS_W-1:0] rs1_phys, rs2_phys, rd_phys, rd_new_phys;

  // -------------------------
  // Instantiate DUT
  // -------------------------
  commit_rename #(
    .ARCH_REGS(ARCH_REGS),
    .PHYS_REGS(PHYS_REGS),
    .ROB_SIZE(ROB_SIZE),
    .ROB_W(ROB_W),
    .PHYS_W(PHYS_W)
  ) dut (
    .clk(clk),
    .rst_n(rst_n),

    .alloc_valid(alloc_valid),
    .alloc_ready(alloc_ready),
    .alloc_uses_rd(alloc_uses_rd),
    .alloc_rd_arch(alloc_rd_arch),
    .alloc_is_branch(alloc_is_branch),
    .alloc_is_load(alloc_is_load),
    .alloc_is_store(alloc_is_store),
    .alloc_pc(alloc_pc),
    .alloc_epoch(alloc_epoch),
    .alloc_rob_idx(alloc_rob_idx),

    .wb_valid(wb_valid),
    .wb_rob_idx(wb_rob_idx),
    .wb_epoch(wb_epoch),

    .commit_valid(commit_valid),
    .commit_ready(commit_ready),

    .commit_uses_rd(commit_uses_rd),
    .commit_rd_arch(commit_rd_arch),
    .commit_pd_new(commit_pd_new),
    .commit_pd_old(commit_pd_old),
    .commit_is_branch(commit_is_branch),
    .commit_is_load(commit_is_load),
    .commit_is_store(commit_is_store),

    .flush_valid(flush_valid),
    .flush_rob_idx(flush_rob_idx),
    .flush_epoch(flush_epoch),

    .rs1_arch(rs1_arch),
    .rs2_arch(rs2_arch),

    .rs1_phys(rs1_phys_dbg),
    .rs2_phys(rs2_phys_dbg),
    .rd_phys(rd_phys_dbg),
    .rd_new_phys(rd_new_phys_dbg)
  );

  always_comb begin
    rs1_phys    = rs1_phys_dbg;
    rs2_phys    = rs2_phys_dbg;
    rd_phys     = rd_phys_dbg;
    rd_new_phys = rd_new_phys_dbg;
  end

  // -------------------------
  // Golden model (TB)
  // -------------------------
  logic [PHYS_W-1:0] golden_rat [ARCH_REGS];
  logic [PHYS_W-1:0] golden_free_q[$];   // FIFO freelist model (p32..p63 plus returned regs >=32)
  logic [PHYS_W-1:0] expect_reuse_q[$];  // regs that should be freed and later reused (>=32)

  typedef struct packed {
    logic              uses_rd;
    logic [4:0]        rd_arch;
    logic [PHYS_W-1:0] pd_new;
    logic [PHYS_W-1:0] pd_old;
    logic [ROB_W-1:0]  rob_idx;
    logic              epoch;
    logic [31:0]       pc;
  } uop_t;

  uop_t inflight_q[$]; // in program order: push at alloc, pop at commit

  uop_t i0, i1, i2, i3, i4;
  int seen_reuse = 0;
  int loops = 0;
  logic [PHYS_W-1:0] target;

  // -------------------------
  // Helpers
  // -------------------------
  task automatic init_signals();
    alloc_valid     = 0;
    alloc_uses_rd   = 0;
    alloc_rd_arch   = '0;
    alloc_is_branch = 0;
    alloc_is_load   = 0;
    alloc_is_store  = 0;
    alloc_pc        = '0;
    alloc_epoch     = 0;

    wb_valid        = 0;
    wb_rob_idx      = '0;
    wb_epoch        = 0;

    commit_ready    = 0;

    flush_valid     = 0;
    flush_rob_idx   = '0;
    flush_epoch     = 0;

    rs1_arch        = 5'd1;  // default probe x1 mapping
    rs2_arch        = 5'd2;  // default probe x2 mapping
  endtask

  task automatic golden_reset();
    int i;
    golden_free_q.delete();
    expect_reuse_q.delete();
    inflight_q.delete();

    for (i = 0; i < ARCH_REGS; i++)
      golden_rat[i] = i[PHYS_W-1:0];

    for (i = 32; i < PHYS_REGS; i++)
      golden_free_q.push_back(i[PHYS_W-1:0]);
  endtask

  task automatic do_reset();
    init_signals();
    rst_n = 0;
    golden_reset();
    repeat (3) @(posedge clk);
    rst_n = 1;
    @(posedge clk);
  endtask

  function automatic logic [PHYS_W-1:0] pop_free();
    logic [PHYS_W-1:0] x;
    if (golden_free_q.size() == 0) $fatal(1, "[TB] Golden freelist empty");
    x = golden_free_q[0];
    golden_free_q.pop_front();
    return x;
  endfunction

  task automatic push_free(input logic [PHYS_W-1:0] pd);
    golden_free_q.push_back(pd);
    expect_reuse_q.push_back(pd); // we expect to see this pd re-allocated later
  endtask

  // One-cycle allocation on negedge to avoid TB/DUT race
  task automatic alloc_inst(
    input  logic        uses_rd,
    input  logic [4:0]  rd_arch,
    input  logic [31:0] pc,
    output uop_t        u
  );
    logic [PHYS_W-1:0] exp_old, exp_new;

    // Compute expected rename result from golden model
    exp_old = golden_rat[rd_arch];
    exp_new = uses_rd ? pop_free() : '0;

    @(negedge clk);
    alloc_valid     = 1'b1;
    alloc_uses_rd   = uses_rd;
    alloc_rd_arch   = rd_arch;
    alloc_is_branch = 1'b0;
    alloc_is_load   = 1'b0;
    alloc_is_store  = 1'b0;
    alloc_pc        = pc;
    alloc_epoch     = alloc_epoch; // keep current

    # 1;
    if (alloc_ready !== 1'b1) begin
      push_free(exp_new);
      $fatal(1, "[TB] alloc_ready=0 when trying to allocate");
    end

    // sample debug rename results during this cycle
    // (if your debug phys ports are too narrow, you'll see truncation here)
    if (uses_rd) begin
      if (rd_phys !== exp_old) $fatal(1, "[TB] Rename pd_old mismatch: exp=%0d got=%0d (rd=x%0d pc=%h)", exp_old, rd_phys, rd_arch, pc);
      if (rd_new_phys !== exp_new) $fatal(1, "[TB] Rename pd_new mismatch: exp=%0d got=%0d (rd=x%0d pc=%h)", exp_new, rd_new_phys, rd_arch, pc);
    end

    // record uop (ROB idx comes from dut output at handshake)
    u.uses_rd = uses_rd;
    u.rd_arch = rd_arch;
    u.pd_old  = exp_old;
    u.pd_new  = exp_new;
    u.rob_idx = alloc_rob_idx;
    u.epoch   = alloc_epoch;
    u.pc      = pc;

    // Update golden RAT after rename
    if (uses_rd) golden_rat[rd_arch] = exp_new;

    inflight_q.push_back(u);

    @(negedge clk);
    alloc_valid = 1'b0;
  endtask

  task automatic wb_done(input logic [ROB_W-1:0] idx, input logic epoch);
    @(negedge clk);
    wb_valid   = 1'b1;
    wb_rob_idx = idx;
    wb_epoch   = epoch;
    @(negedge clk);
    wb_valid   = 1'b0;
  endtask

  task automatic commit_one();
    uop_t u;
    int watchdog = 0;

    if (inflight_q.size() == 0) $fatal(1, "[TB] commit_one: inflight empty");
    u = inflight_q[0];

    // wait for commit_valid
    while (!commit_valid) begin
      @(posedge clk);
      watchdog++;
      if (watchdog > 200) $fatal(1, "[TB] Timeout waiting commit_valid");
    end

    // accept commit
    @(negedge clk);
    commit_ready = 1'b1;
    @(negedge clk);
    commit_ready = 1'b0;

    // Check commit fields (architectural retirement order)
    if (commit_uses_rd !== u.uses_rd) $fatal(1, "[TB] commit_uses_rd mismatch");
    if (u.uses_rd) begin
      if (commit_rd_arch !== u.rd_arch) $fatal(1, "[TB] commit_rd_arch mismatch exp=x%0d got=x%0d pc=%h", u.rd_arch, commit_rd_arch, u.pc);
      if (commit_pd_new  !== u.pd_new)  $fatal(1, "[TB] commit_pd_new mismatch exp=%0d got=%0d pc=%h", u.pd_new, commit_pd_new, u.pc);
      if (commit_pd_old  !== u.pd_old)  $fatal(1, "[TB] commit_pd_old mismatch exp=%0d got=%0d pc=%h", u.pd_old, commit_pd_old, u.pc);

      // Golden: on commit, free pd_old (if >=32)
      push_free(u.pd_old);
    end

    inflight_q.pop_front();
  endtask

  // -------------------------
  // Extra TB helpers / tests
  // -------------------------

  // Drive an allocation attempt and EXPECT alloc_ready=0 (no handshake should occur).
  task automatic alloc_expect_stall(
    input logic        uses_rd,
    input logic [4:0]  rd_arch,
    input logic [31:0] pc
  );
    int free_sz_before;
    free_sz_before = golden_free_q.size();

    @(negedge clk);
    alloc_valid     = 1'b1;
    alloc_uses_rd   = uses_rd;
    alloc_rd_arch   = rd_arch;
    alloc_is_branch = 1'b0;
    alloc_is_load   = 1'b0;
    alloc_is_store  = 1'b0;
    alloc_pc        = pc;
    alloc_epoch     = alloc_epoch;

    // Give the DUT a delta to resolve ready/outputs.
    #1;
    if (alloc_ready !== 1'b0) begin
      $fatal(1, "[TB] Expected alloc_ready=0 (stall) but got alloc_ready=1 at pc=%h rd=x%0d", pc, rd_arch);
    end
    // Golden model must not change on a stall
    if (golden_free_q.size() !== free_sz_before) begin
      $fatal(1, "[TB] Golden freelist changed during a supposed stall");
    end

    @(negedge clk);
    alloc_valid = 1'b0;
  endtask

  // Fill the ROB (or other alloc-side resource) and ensure alloc_ready deasserts.
  // This is a practical substitute for "freelist empty" when ROB_SIZE < (#free phys regs).
  task automatic test_rob_full_stall();
    uop_t tmp;
    int i;

    $display("=== TEST B: Fill ROB and ensure alloc stalls when full ===");

    // Fill to ROB_SIZE inflight uops without writeback/commit.
    for (i = 0; i < ROB_SIZE; i++) begin
      alloc_inst(1'b1, 5'd1, 32'h2000 + 4*i, tmp);
    end

    // Next allocate should stall (alloc_ready=0). If your DUT also gates on freelist, this still holds.
    alloc_expect_stall(1'b1, 5'd2, 32'h3000);

    // Now retire one uop to create space and ensure alloc resumes.
    wb_done(inflight_q[0].rob_idx, inflight_q[0].epoch);
    commit_one();

    // Should be able to allocate again now.
    alloc_inst(1'b1, 5'd2, 32'h3004, tmp);

    // Clean up: retire everything we left inflight to avoid polluting later tests.
    while (inflight_q.size() != 0) begin
      wb_done(inflight_q[0].rob_idx, inflight_q[0].epoch);
      commit_one();
    end
  endtask

  // Sanity: an instruction with no destination must not consume a physical register.
  task automatic test_no_rd_does_not_allocate();
    uop_t u;
    int free_before, free_after;

    $display("=== TEST C: uses_rd=0 does not pop freelist ===");

    free_before = golden_free_q.size();
    alloc_inst(1'b0, 5'd0, 32'h4000, u);
    free_after  = golden_free_q.size();

    if (free_after !== free_before) begin
      $fatal(1, "[TB] uses_rd=0 changed freelist size: before=%0d after=%0d", free_before, free_after);
    end

    // If it allocates into ROB, still needs commit path; complete it.
    wb_done(u.rob_idx, u.epoch);
    commit_one();
  endtask


  // -------------------------
  // Cycle-by-cycle display
  // -------------------------
  always @(posedge clk) begin
    if (rst_n & alloc_valid) begin
      $display("[C%0t] alloc_v=%0d rdy=%0d rd=x%0d old=%0d new=%0d | rs1=x%0d->p%0d rs2=x%0d->p%0d | commit_v=%0d",
        $time, alloc_valid, alloc_ready, alloc_rd_arch, rd_phys, rd_new_phys,
        rs1_arch, rs1_phys, rs2_arch, rs2_phys,
        commit_valid
      );
    end
    else if (rst_n & commit_valid & commit_ready) begin
      $display("[C%0t] committing instn | rs1=x%0d->p%0d rs2=x%0d->p%0d | commit_v=%0d rd=x%0d old=%0d new=%0d",
        $time,
        rs1_arch, rs1_phys, rs2_arch, rs2_phys,
        commit_valid,
        commit_rd_arch, commit_pd_old, commit_pd_new
      );
    end
  end

  // -------------------------
  // Main tests
  // -------------------------
  initial begin
    do_reset();

    // If debug phys ports are only 5 bits, they cannot show p32..p63 correctly.
    // Warn once if we detect truncation (rd_new_phys should become >=32 quickly).
    @(negedge clk);

    // ---- TEST A: WAW + RAW hazard case and correct commit freeing/reuse ----
    // I0: x1 = ...
    // I1: x1 = ...
    // I2: r = x1  (we check mapping by probing rs1_arch=x1 at rename time)

    rs1_arch = 5'd1; // probe x1 mapping
    rs2_arch = 5'd2; // probe x2 mapping

    $display("=== TEST A: WAW then probe RAW mapping ===");
    alloc_inst(1'b1, 5'd1, 32'h1000, i0); // expects old=p1 new=p32
    alloc_inst(1'b1, 5'd1, 32'h1004, i1); // expects old=p32 new=p33
    // After I1 rename, RAT[x1] should be p33, so rs1_phys should show p33 when probing x1
    @(negedge clk);
    if (rs1_phys !== golden_rat[1]) $fatal(1, "[TB] RAT probe mismatch after WAW: exp p%0d got p%0d", golden_rat[1], rs1_phys);

    // Mark writebacks out of order to ensure commit is still in order
    wb_done(i1.rob_idx, i1.epoch);
    wb_done(i0.rob_idx, i0.epoch);

    // Commit in order (I0 then I1)
    commit_one(); // commits I0 -> frees p1? (ignored because <32)
    commit_one(); // commits I1 -> frees p32 (should reappear later)

    // Now allocate a few more to eventually observe p32 reused
    $display("=== Alloc more to observe freed reg reuse ===");
    alloc_inst(1'b1, 5'd2, 32'h1010, i2); // x2 writer
    alloc_inst(1'b1, 5'd3, 32'h1014, i3); // x3 writer
    alloc_inst(1'b1, 5'd4, 32'h1018, i4); // x4 writer

    // complete + commit these
    wb_done(i2.rob_idx, i2.epoch);
    wb_done(i3.rob_idx, i3.epoch);
    wb_done(i4.rob_idx, i4.epoch);
    commit_one();
    commit_one();
    commit_one();

    // Check that a freed reg (p32) is eventually reallocated as a future pd_new.
    // We track expected_reuse_q; simplest check: after some allocs, see one of them appear.
    // Allocate until we see a re-used pd (bounded loop).
    if (expect_reuse_q.size() > 0) target = expect_reuse_q[0];

    while (!seen_reuse && loops < 40) begin
      uop_t t;
      alloc_inst(1'b1, 5'd5, 32'h2000 + loops*4, t);
      if (t.pd_new == target) begin
        $display("[TB] Observed freed pd_old p%0d re-allocated as pd_new ✅", target);
        seen_reuse = 1;
      end
      // make it commit quickly
      wb_done(t.rob_idx, t.epoch);
      commit_one();
      loops++;
    end

    if (!seen_reuse) begin
      $fatal(1, "[TB] Did not observe freed pd_old p%0d being reused within bound. Either freelist not freeing or FIFO order differs.", target);
    end

    // ---- TEST B: Fill ROB and ensure alloc stalls when full ----
    test_rob_full_stall();
    // ---- TEST C: uses_rd=0 does not consume physical register ----
    test_no_rd_does_not_allocate();

    $display("[TB] ALL COMMIT+RENAME TESTS PASS ✅");
    $finish;
  end

endmodule
